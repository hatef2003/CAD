`timescale 1ps/1ps
module eight_bit_adder( input [11:0] a , b , output [11:0] result);
    assign result = a + b ;
endmodule