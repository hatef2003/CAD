module Xor (input a , b , output o);
 c2 cell1(0,1,1,0,a,b,a,b,o);
endmodule